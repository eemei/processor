library verilog;
use verilog.vl_types.all;
entity addTB is
end addTB;

module register8bitTB ();
  wire [7:0] Q; 
 reg [7:0] D;
 reg load, Clock, Reset;

 
initial 
begin 
Clock = 0;
Reset = 0;
load = 0;
D= 0;
#7 Reset =1; load =1;
#4 D = 8'b00000110;
#4 D = 8'b11001011;
#4 D = 8'b11011;
#20 $finish;
end

always @(Q)begin
$display("OUTPUT IR= %b", Q);
end

always #1 Clock = ~Clock;

register8bit  #(.SIZE(8))regTB(Q,D,load,Clock,Reset);
//register8bit  #(.SIZE(5))regTB_5(IR,D,IRload,Clock,Reset);
 
endmodule

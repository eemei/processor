library verilog;
use verilog.vl_types.all;
entity CUtb is
end CUtb;

library verilog;
use verilog.vl_types.all;
entity IRregTB is
end IRregTB;

library verilog;
use verilog.vl_types.all;
entity RAMtb is
end RAMtb;

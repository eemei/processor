library verilog;
use verilog.vl_types.all;
entity Aregistertb is
end Aregistertb;

library verilog;
use verilog.vl_types.all;
entity BarrelTB is
end BarrelTB;
